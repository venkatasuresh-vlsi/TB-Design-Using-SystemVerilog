module matrix_mul(
     input [3:0] a[3:0][3:0],
     input [3:0] b[3:0][3:0],
	 output [15:0] y[3:0][3:0]
	 );
	 assign y[0][0] =
	    (a[0][0] * b[0][0]) +
		(a[0][1] * b[1][0]) +
		(a[0][2] * b[2][0]) +
		(a[0][3] * b[3][0]) ;
	 assign y[0][1] =
		(a[0][0] * b[0][1]) +
		(a[0][1] * b[1][1]) +
		(a[0][2] * b[2][1]) +
		(a[0][3] * b[3][1]) ;
	 assign y[0][2] =
		(a[0][0] * b[0][2]) +
		(a[0][1] * b[1][2]) +
		(a[0][2] * b[2][2]) +
		(a[0][3] * b[3][2]) ;
	 assign y[0][3] =
		(a[0][0] * b[0][3]) +
		(a[0][1] * b[1][3]) +
		(a[0][2] * b[2][3]) +
		(a[0][3] * b[3][3]) ;
	 assign y[1][0] =
		(a[1][0] * b[0][0]) +
		(a[1][1] * b[1][0]) +
		(a[1][2] * b[2][0]) +
		(a[1][3] * b[3][0]) ;
	 assign y[1][1] =
		(a[1][0] * b[0][1]) +
		(a[1][1] * b[1][1]) +
		(a[1][2] * b[2][1]) +
		(a[1][3] * b[3][1]) ;
	 assign y[1][2] =
		(a[1][0] * b[0][2]) +
		(a[1][1] * b[1][2]) +
		(a[1][2] * b[2][2]) +
		(a[1][3] * b[3][2]) ;
	 assign y[1][3] =
		(a[1][0] * b[0][3]) +
		(a[1][1] * b[1][3]) +
		(a[1][2] * b[2][3]) +
		(a[1][3] * b[3][3]) ;
	 assign y[2][0] =
		(a[2][0] * b[0][0]) +
		(a[2][1] * b[1][0]) +
		(a[2][2] * b[2][0]) +
		(a[2][3] * b[3][0]) ;
	 assign y[2][1] =
		(a[2][0] * b[0][1]) +
		(a[2][1] * b[1][1]) +
		(a[2][2] * b[2][1]) +
		(a[2][3] * b[3][1]) ;
	 assign y[2][2] =
		(a[2][0] * b[0][2]) +
		(a[2][1] * b[1][2]) +
		(a[2][2] * b[2][2]) +
		(a[2][3] * b[3][2]) ;
	 assign y[2][3] =
		(a[2][0] * b[0][3]) +
		(a[2][1] * b[1][3]) +
		(a[2][2] * b[2][3]) +
		(a[2][3] * b[3][3]) ;
	 assign y[3][0] =
		(a[3][0] * b[0][0]) +
		(a[3][1] * b[1][0]) +
		(a[3][2] * b[2][0]) +
		(a[3][3] * b[3][0]) ;
	 assign y[3][1] =
		(a[3][0] * b[0][1]) +
		(a[3][1] * b[1][1]) +
		(a[3][2] * b[2][1]) +
		(a[3][3] * b[3][1]) ;
	 assign y[3][2] =
		(a[3][0] * b[0][2]) +
		(a[3][1] * b[1][2]) +
		(a[3][2] * b[2][2]) +
		(a[3][3] * b[3][2]) ;
	 assign y[3][3] =
		(a[3][0] * b[0][3]) +
		(a[3][1] * b[1][3]) +
		(a[3][2] * b[2][3]) +
		(a[3][3] * b[3][3]) ;
    
	endmodule