class mux_connections;
     rand bit [3:0] a;
     rand bit [3:0] b;
	 rand bit sel;
	      bit [3:0] y;
	endclass